class transaction;
    rand bit cnt;
        bit[7:0] din;
        bit wr;
        bit rd;
        bit full;
        bit empty;
        bit[7:0] dut;

        constraint dist{
endclass
