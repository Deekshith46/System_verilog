interface dff();
    logic din;
    logic dout;
    logic clk;
    logic rst;
endinterface
