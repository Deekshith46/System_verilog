class transaction;

    rand bit din;
    bit dout;

    function transaction copy();
        copy = new();
        copy.din = this.din;
        copy.dout = this.dout;
    endfunction

    function void display(input string tag);
        $display("[%0s]: DIN : %0b DOUT : %0b",tag,din,dout);
    endfunction
    
endclass
